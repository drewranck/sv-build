
`ifndef sv_build_example_includes__svh
`define sv_build_example_includes__svh

`include "sv_build_example_srl_defines.svh"

`endif
